--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package text_package is
	
	type point_2d is
	record
		x : integer;
		y : integer;
	end record;

	type type_text_lineDebug is
	record
		debugDraw: std_logic_vector(39 downto 0);
	end record;

--	type type_characterMap is array (character) of std_logic_vector(7 downto 0);
--	constant ascii_address_xref : type_characterMap := (
--		-- Char => Addr	-- Decimal : Hex
--		character'val(16#00#) => "00000000",	-- NULL : 0 : x00
--		character'val(16#01#) => "00000001",	--  : 1 : x01
--		character'val(16#02#) => "00000010",	--  : 2 : x02
--		character'val(16#03#) => "00000011",	--  : 3 : x03
--		character'val(16#04#) => "00000100",	--  : 4 : x04
--		character'val(16#05#) => "00000101",	--  : 5 : x05
--		character'val(16#06#) => "00000110",	--  : 6 : x06
--		character'val(16#07#) => "00000111",	--  : 7 : x07
--		character'val(16#08#) => "00001000",	--  : 8 : x08
--		character'val(16#09#) => "00001001",	-- HT Tab : 9 : x09
--		character'val(16#0a#) => "00001010",	-- LF : 10 : x0a
--		character'val(16#0b#) => "00001011",	--  : 11 : x0b
--		character'val(16#0c#) => "00001100",	--  : 12 : x0c
--		character'val(16#0d#) => "00001101",	-- CR : 13 : x0d
--		character'val(16#0e#) => "00001110",	--  : 14 : x0e
--		character'val(16#0f#) => "00001111",	--  : 15 : x0f
--		character'val(16#10#) => "00010000",	--  : 16 : x10
--		character'val(16#11#) => "00010001",	--  : 17 : x11
--		character'val(16#12#) => "00010010",	--  : 18 : x12
--		character'val(16#13#) => "00010011",	--  : 19 : x13
--		character'val(16#14#) => "00010100",	--  : 20 : x14
--		character'val(16#15#) => "00010101",	--  : 21 : x15
--		character'val(16#16#) => "00010110",	--  : 22 : x16
--		character'val(16#17#) => "00010111",	--  : 23 : x17
--		character'val(16#18#) => "00011000",	--  : 24 : x18
--		character'val(16#19#) => "00011001",	--  : 25 : x19
--		character'val(16#1a#) => "00011010",	--  : 26 : x1a
--		character'val(16#1b#) => "00011011",	--  : 27 : x1b
--		character'val(16#1c#) => "00011100",	--  : 28 : x1c
--		character'val(16#1d#) => "00011101",	--  : 29 : x1d
--		character'val(16#1e#) => "00011110",	--  : 30 : x1e
--		character'val(16#1f#) => "00011111",	--  : 31 : x1f
--		character'val(16#20#) => "00100000",	-- SP Space : 32 : x20
--		character'val(16#21#) => "00100001",	-- ! : 33 : x21
--		character'val(16#22#) => "00100010",	-- " : 34 : x22
--		character'val(16#23#) => "00100011",	-- # : 35 : x23
--		character'val(16#24#) => "00100100",	-- $ : 36 : x24
--		character'val(16#25#) => "00100101",	-- % : 37 : x25
--		character'val(16#26#) => "00100110",	-- & : 38 : x26
--		character'val(16#27#) => "00100111",	-- ' : 39 : x27
--		character'val(16#28#) => "00101000",	-- ( : 40 : x28
--		character'val(16#29#) => "00101001",	-- ) : 41 : x29
--		character'val(16#2a#) => "00101010",	-- * : 42 : x2a
--		character'val(16#2b#) => "00101011",	-- + : 43 : x2b
--		character'val(16#2c#) => "00101100",	-- , : 44 : x2c
--		character'val(16#2d#) => "00101101",	-- - : 45 : x2d
--		character'val(16#2e#) => "00101110",	-- . : 46 : x2e
--		character'val(16#2f#) => "00101111",	-- / : 47 : x2f
--		character'val(16#30#) => "00110000",	-- 0 : 48 : x30
--		character'val(16#31#) => "00110001",	-- 1 : 49 : x31
--		character'val(16#32#) => "00110010",	-- 2 : 50 : x32
--		character'val(16#33#) => "00110011",	-- 3 : 51 : x33
--		character'val(16#34#) => "00110100",	-- 4 : 52 : x34
--		character'val(16#35#) => "00110101",	-- 5 : 53 : x35
--		character'val(16#36#) => "00110110",	-- 6 : 54 : x36
--		character'val(16#37#) => "00110111",	-- 7 : 55 : x37
--		character'val(16#38#) => "00111000",	-- 8 : 56 : x38
--		character'val(16#39#) => "00111001",	-- 9 : 57 : x39
--		character'val(16#3a#) => "00111010",	-- : : 58 : x3a
--		character'val(16#3b#) => "00111011",	-- ; : 59 : x3b
--		character'val(16#3c#) => "00111100",	-- < : 60 : x3c
--		character'val(16#3d#) => "00111101",	-- = : 61 : x3d
--		character'val(16#3e#) => "00111110",	-- > : 62 : x3e
--		character'val(16#3f#) => "00111111",	-- ? : 63 : x3f
--		character'val(16#40#) => "01000000",	-- @ : 64 : x40
--		character'val(16#41#) => "01000001",	-- A : 65 : x41
--		character'val(16#42#) => "01000010",	-- B : 66 : x42
--		character'val(16#43#) => "01000011",	-- C : 67 : x43
--		character'val(16#44#) => "01000100",	-- D : 68 : x44
--		character'val(16#45#) => "01000101",	-- E : 69 : x45
--		character'val(16#46#) => "01000110",	-- F : 70 : x46
--		character'val(16#47#) => "01000111",	-- G : 71 : x47
--		character'val(16#48#) => "01001000",	-- H : 72 : x48
--		character'val(16#49#) => "01001001",	-- I : 73 : x49
--		character'val(16#4a#) => "01001010",	-- J : 74 : x4a
--		character'val(16#4b#) => "01001011",	-- K : 75 : x4b
--		character'val(16#4c#) => "01001100",	-- L : 76 : x4c
--		character'val(16#4d#) => "01001101",	-- M : 77 : x4d
--		character'val(16#4e#) => "01001110",	-- N : 78 : x4e
--		character'val(16#4f#) => "01001111",	-- O : 79 : x4f
--		character'val(16#50#) => "01010000",	-- P : 80 : x50
--		character'val(16#51#) => "01010001",	-- Q : 81 : x51
--		character'val(16#52#) => "01010010",	-- R : 82 : x52
--		character'val(16#53#) => "01010011",	-- S : 83 : x53
--		character'val(16#54#) => "01010100",	-- T : 84 : x54
--		character'val(16#55#) => "01010101",	-- U : 85 : x55
--		character'val(16#56#) => "01010110",	-- V : 86 : x56
--		character'val(16#57#) => "01010111",	-- W : 87 : x57
--		character'val(16#58#) => "01011000",	-- X : 88 : x58
--		character'val(16#59#) => "01011001",	-- Y : 89 : x59
--		character'val(16#5a#) => "01011010",	-- Z : 90 : x5a
--		character'val(16#5b#) => "01011011",	-- [ : 91 : x5b
--		character'val(16#5c#) => "01011100",	-- \ : 92 : x5c
--		character'val(16#5d#) => "01011101",	-- ] : 93 : x5d
--		character'val(16#5e#) => "01011110",	-- ^ : 94 : x5e
--		character'val(16#5f#) => "01011111",	-- _ : 95 : x5f
--		character'val(16#60#) => "01100000",	-- ` : 96 : x60
--		character'val(16#61#) => "01100001",	-- a : 97 : x61
--		character'val(16#62#) => "01100010",	-- b : 98 : x62
--		character'val(16#63#) => "01100011",	-- c : 99 : x63
--		character'val(16#64#) => "01100100",	-- d : 100 : x64
--		character'val(16#65#) => "01100101",	-- e : 101 : x65
--		character'val(16#66#) => "01100110",	-- f : 102 : x66
--		character'val(16#67#) => "01100111",	-- g : 103 : x67
--		character'val(16#68#) => "01101000",	-- h : 104 : x68
--		character'val(16#69#) => "01101001",	-- i : 105 : x69
--		character'val(16#6a#) => "01101010",	-- j : 106 : x6a
--		character'val(16#6b#) => "01101011",	-- k : 107 : x6b
--		character'val(16#6c#) => "01101100",	-- l : 108 : x6c
--		character'val(16#6d#) => "01101101",	-- m : 109 : x6d
--		character'val(16#6e#) => "01101110",	-- n : 110 : x6e
--		character'val(16#6f#) => "01101111",	-- o : 111 : x6f
--		character'val(16#70#) => "01110000",	-- p : 112 : x70
--		character'val(16#71#) => "01110001",	-- q : 113 : x71
--		character'val(16#72#) => "01110010",	-- r : 114 : x72
--		character'val(16#73#) => "01110011",	-- s : 115 : x73
--		character'val(16#74#) => "01110100",	-- t : 116 : x74
--		character'val(16#75#) => "01110101",	-- u : 117 : x75
--		character'val(16#76#) => "01110110",	-- v : 118 : x76
--		character'val(16#77#) => "01110111",	-- w : 119 : x77
--		character'val(16#78#) => "01111000",	-- x : 120 : x78
--		character'val(16#79#) => "01111001",	-- y : 121 : x79
--		character'val(16#7a#) => "01111010",	-- z : 122 : x7a
--		character'val(16#7b#) => "01111011",	-- { : 123 : x7b
--		character'val(16#7c#) => "01111100",	-- | : 124 : x7c
--		character'val(16#7d#) => "01111101",	-- } : 125 : x7d
--		character'val(16#7e#) => "01111110",	-- ~ : 126 : x7e
--		character'val(16#7f#) => "01111111",	-- DEL : 127 : x7f
--		character'val(16#80#) => "10000000",	-- � : 128 : x80
--		character'val(16#81#) => "10000001",	-- HOP	High Octet Preset : 129 : x81
--		character'val(16#82#) => "10000010",	-- � : 130 : x82
--		character'val(16#83#) => "10000011",	-- � : 131 : x83
--		character'val(16#84#) => "10000100",	-- � : 132 : x84
--		character'val(16#85#) => "10000101",	-- � : 133 : x85
--		character'val(16#86#) => "10000110",	-- � : 134 : x86
--		character'val(16#87#) => "10000111",	-- � : 135 : x87
--		character'val(16#88#) => "10001000",	-- � : 136 : x88
--		character'val(16#89#) => "10001001",	-- � : 137 : x89
--		character'val(16#8a#) => "10001010",	-- � : 138 : x8a
--		character'val(16#8b#) => "10001011",	-- � : 139 : x8b
--		character'val(16#8c#) => "10001100",	-- � : 140 : x8c
--		character'val(16#8d#) => "10001101",	-- � : 141 : x8d
--		character'val(16#8e#) => "10001110",	-- � : 142 : x8e
--		character'val(16#8f#) => "10001111",	-- SS3	Single Shift 3 : 143 : x8f
--		character'val(16#90#) => "10010000",	-- DCS	Device Control String : 144 : x90
--		character'val(16#91#) => "10010001",	-- ' : 145 : x91
--		character'val(16#92#) => "10010010",	-- ' : 146 : x92
--		character'val(16#93#) => "10010011",	-- " : 147 : x93
--		character'val(16#94#) => "10010100",	-- " : 148 : x94
--		character'val(16#95#) => "10010101",	-- � : 149 : x95
--		character'val(16#96#) => "10010110",	-- - : 150 : x96
--		character'val(16#97#) => "10010111",	-- - : 151 : x97
--		character'val(16#98#) => "10011000",	-- � : 152 : x98
--		character'val(16#99#) => "10011001",	-- � : 153 : x99
--		character'val(16#9a#) => "10011010",	-- � : 154 : x9a
--		character'val(16#9b#) => "10011011",	-- � : 155 : x9b
--		character'val(16#9c#) => "10011100",	-- � : 156 : x9c
--		character'val(16#9d#) => "10011101",	-- OSC	Operating System Command : 157 : x9d
--		character'val(16#9e#) => "10011110",	-- � : 158 : x9e
--		character'val(16#9f#) => "10011111",	-- � : 159 : x9f
--		character'val(16#a0#) => "10100000",	-- NBSP Space : 160 : xa0
--		character'val(16#a1#) => "10100001",	-- � : 161 : xa1
--		character'val(16#a2#) => "10100010",	-- � : 162 : xa2
--		character'val(16#a3#) => "10100011",	-- � : 163 : xa3
--		character'val(16#a4#) => "10100100",	-- � : 164 : xa4
--		character'val(16#a5#) => "10100101",	-- � : 165 : xa5
--		character'val(16#a6#) => "10100110",	-- � : 166 : xa6
--		character'val(16#a7#) => "10100111",	-- � : 167 : xa7
--		character'val(16#a8#) => "10101000",	-- � : 168 : xa8
--		character'val(16#a9#) => "10101001",	-- � : 169 : xa9
--		character'val(16#aa#) => "10101010",	-- � : 170 : xaa
--		character'val(16#ab#) => "10101011",	-- � : 171 : xab
--		character'val(16#ac#) => "10101100",	-- � : 172 : xac
--		character'val(16#ad#) => "10101101",	-- � : 173 : xad
--		character'val(16#ae#) => "10101110",	-- � : 174 : xae
--		character'val(16#af#) => "10101111",	-- � : 175 : xaf
--		character'val(16#b0#) => "10110000",	-- � : 176 : xb0
--		character'val(16#b1#) => "10110001",	-- � : 177 : xb1
--		character'val(16#b2#) => "10110010",	-- � : 178 : xb2
--		character'val(16#b3#) => "10110011",	-- � : 179 : xb3
--		character'val(16#b4#) => "10110100",	-- � : 180 : xb4
--		character'val(16#b5#) => "10110101",	-- � : 181 : xb5
--		character'val(16#b6#) => "10110110",	-- � : 182 : xb6
--		character'val(16#b7#) => "10110111",	-- � : 183 : xb7
--		character'val(16#b8#) => "10111000",	-- � : 184 : xb8
--		character'val(16#b9#) => "10111001",	-- � : 185 : xb9
--		character'val(16#ba#) => "10111010",	-- � : 186 : xba
--		character'val(16#bb#) => "10111011",	-- � : 187 : xbb
--		character'val(16#bc#) => "10111100",	-- � : 188 : xbc
--		character'val(16#bd#) => "10111101",	-- � : 189 : xbd
--		character'val(16#be#) => "10111110",	-- � : 190 : xbe
--		character'val(16#bf#) => "10111111",	-- � : 191 : xbf
--		character'val(16#c0#) => "11000000",	-- � : 192 : xc0
--		character'val(16#c1#) => "11000001",	-- � : 193 : xc1
--		character'val(16#c2#) => "11000010",	-- � : 194 : xc2
--		character'val(16#c3#) => "11000011",	-- � : 195 : xc3
--		character'val(16#c4#) => "11000100",	-- � : 196 : xc4
--		character'val(16#c5#) => "11000101",	-- � : 197 : xc5
--		character'val(16#c6#) => "11000110",	-- � : 198 : xc6
--		character'val(16#c7#) => "11000111",	-- � : 199 : xc7
--		character'val(16#c8#) => "11001000",	-- � : 200 : xc8
--		character'val(16#c9#) => "11001001",	-- � : 201 : xc9
--		character'val(16#ca#) => "11001010",	-- � : 202 : xca
--		character'val(16#cb#) => "11001011",	-- � : 203 : xcb
--		character'val(16#cc#) => "11001100",	-- � : 204 : xcc
--		character'val(16#cd#) => "11001101",	-- � : 205 : xcd
--		character'val(16#ce#) => "11001110",	-- � : 206 : xce
--		character'val(16#cf#) => "11001111",	-- � : 207 : xcf
--		character'val(16#d0#) => "11010000",	-- � : 208 : xd0
--		character'val(16#d1#) => "11010001",	-- � : 209 : xd1
--		character'val(16#d2#) => "11010010",	-- � : 210 : xd2
--		character'val(16#d3#) => "11010011",	-- � : 211 : xd3
--		character'val(16#d4#) => "11010100",	-- � : 212 : xd4
--		character'val(16#d5#) => "11010101",	-- � : 213 : xd5
--		character'val(16#d6#) => "11010110",	-- � : 214 : xd6
--		character'val(16#d7#) => "11010111",	-- � : 215 : xd7
--		character'val(16#d8#) => "11011000",	-- � : 216 : xd8
--		character'val(16#d9#) => "11011001",	-- � : 217 : xd9
--		character'val(16#da#) => "11011010",	-- � : 218 : xda
--		character'val(16#db#) => "11011011",	-- � : 219 : xdb
--		character'val(16#dc#) => "11011100",	-- � : 220 : xdc
--		character'val(16#dd#) => "11011101",	-- � : 221 : xdd
--		character'val(16#de#) => "11011110",	-- � : 222 : xde
--		character'val(16#df#) => "11011111",	-- � : 223 : xdf
--		character'val(16#e0#) => "11100000",	-- � : 224 : xe0
--		character'val(16#e1#) => "11100001",	-- � : 225 : xe1
--		character'val(16#e2#) => "11100010",	-- � : 226 : xe2
--		character'val(16#e3#) => "11100011",	-- � : 227 : xe3
--		character'val(16#e4#) => "11100100",	-- � : 228 : xe4
--		character'val(16#e5#) => "11100101",	-- � : 229 : xe5
--		character'val(16#e6#) => "11100110",	-- � : 230 : xe6
--		character'val(16#e7#) => "11100111",	-- � : 231 : xe7
--		character'val(16#e8#) => "11101000",	-- � : 232 : xe8
--		character'val(16#e9#) => "11101001",	-- � : 233 : xe9
--		character'val(16#ea#) => "11101010",	-- � : 234 : xea
--		character'val(16#eb#) => "11101011",	-- � : 235 : xeb
--		character'val(16#ec#) => "11101100",	-- � : 236 : xec
--		character'val(16#ed#) => "11101101",	-- � : 237 : xed
--		character'val(16#ee#) => "11101110",	-- � : 238 : xee
--		character'val(16#ef#) => "11101111",	-- � : 239 : xef
--		character'val(16#f0#) => "11110000",	-- � : 240 : xf0
--		character'val(16#f1#) => "11110001",	-- � : 241 : xf1
--		character'val(16#f2#) => "11110010",	-- � : 242 : xf2
--		character'val(16#f3#) => "11110011",	-- � : 243 : xf3
--		character'val(16#f4#) => "11110100",	-- � : 244 : xf4
--		character'val(16#f5#) => "11110101",	-- � : 245 : xf5
--		character'val(16#f6#) => "11110110",	-- � : 246 : xf6
--		character'val(16#f7#) => "11110111",	-- � : 247 : xf7
--		character'val(16#f8#) => "11111000",	-- � : 248 : xf8
--		character'val(16#f9#) => "11111001",	-- � : 249 : xf9
--		character'val(16#fa#) => "11111010",	-- � : 250 : xfa
--		character'val(16#fb#) => "11111011",	-- � : 251 : xfb
--		character'val(16#fc#) => "11111100",	-- � : 252 : xfc
--		character'val(16#fd#) => "11111101",	-- � : 253 : xfd
--		character'val(16#fe#) => "11111110",	-- � : 254 : xfe
--		character'val(16#ff#) => "11111111"		-- � : 255 : xff
--	);

end text_package;

package body text_package is

 
end text_package;
